library verilog;
use verilog.vl_types.all;
entity adder64_vlg_vec_tst is
end adder64_vlg_vec_tst;
