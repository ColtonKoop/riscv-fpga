module arithmetic_unit()

endmodule 